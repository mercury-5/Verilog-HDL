module and_gt (y, a, b);
    
    input a, b;
    output y;

and A1(y, a, b);

endmodule